`timescale 1ns/1ps

package test_regs_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  import gr_reg_pkg::*;
  
  `include "sv/register/test_reg_model.sv"
   
  //`include "sv/test_seq.sv"
endpackage
