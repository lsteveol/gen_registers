//===================================================================
//
// Copyright (C) Wavious 2019 - All Rights Reserved
//
// Unauthorized copying of this file, via any medium is strictly prohibited
//
// Created by sbridges on November/11/2019 at 13:18:06
//
// wav_reg_model_lss_no_reg_test.svh
//
//===================================================================






